� �   @������������������������������������������                                     �������������������������������������������                                     ��������������������������������������������                                    ��������������������������������������������                                    ���������������������   �������������������                                    ������������������������������������������                                    ��������������������������Ј����������������                                    ���������������������������Ј����������������                                   ��������������������������������������������                                   ��������������������������������������������                                   ��������������������ݍ������Ј��������������                                   ������������������ݍ�������Ј���������������                                   ������������������ݍ�������������������������                                  ������������������ݍ��ݍ���������������������                                  ��������������������ƍ����������������������                                  �����������������݀��`���������������������                                  �������������������`��n���������������������                                 ������������������ f��o�����Ј����������������                                 ����������������������������������������������                                 �������������������������������������� ������                                 ������������������ؠ��o�nf����Ј���������������                                 �������������������n��f��f����Ј���������������                                �������������������n�Fn��f�����Ј��������������                                �������������������������f`����܍��������������                                ��������������������L���f`�������������������                                ����������������������N��f ������Ј�������������                                ������������������������``������Ј��������������                               �����������������������`f`���������������������                               ���������������������� fff�������������������                               ����������������������ffnf������Ј������������                               ����������������������fn��`-�������������������                               �������������������݈������f#  ������������������                              �����������������݆�"f����fn#.�������������������                              ����������������݆��2�������'.�����Ј������������                              �����������������n��r�������'2������������������                              ��������������������r�������'r���m����������������                             ��������������������r�������'r���ਈ���������������                             �������������������r�������#r���� ���   ��������                             ����        �����r�������#r���h�����   �������                             ������������Ѐ����3.������#r���`������  ��������                             ������������Ѐ����3.������#3.n�`������  ���������                            ����������������b32������'3 n�`������  ���������                            �����������������ws.�f��#ww&n��������  ��������                            ������������������#www2""7wwwrn�������� ��������                            ������������������'wwwwwwwwwwsn�������� ���������                            ����������������.��7wwwwwwwwwww&�������� ����������                           ����������������n�b7wwwwwwwwwww2�������� ����������                           ������������������#7wwwwwwwwwww3.�`������ ���������                           ������������������37wwwwwwwwwws3&�`�����������������                           ������������������33wwwwwwwwwws3&``������������������                          ������������������237www3337ws33&n������������������                          �����������������33333333333332fnf`�����������������                          ���������������nf#333337ww#333 f������������������                          ���������������h f#3"3wwwws2"3
�������������������                          ���������������n�f337wwwwws33 `��������������������                         ���������������fn�f33wwwwwwws3��������������������                         ���������������fn��`337wwwwwws3`�������������������                         ���������������fn�f`'w"�wwwww33�������������������                         ���������������ff�f'wwz#wws2"w�`�����������������                         ���������������fn`
����z#3'���� ��������������������                        ���������������n�� ���zr2��p a`���������������������                        ���������������n�`"" ���*�""  �������������������                        ����������������n�f"""" p """" ` �������������������                        ����������������n��"""""  """""" 0���������������������                       ���������������f���"""""""""""" 0������� ��������������                       ���������������n��� """"""""""2������ ��������������                       ����������������n� ff`"""""""""   ������ �������������                       ����������������n��f"""""""""
fff������ ��������������                       �����������������  """""""" �n�f`������ ���������������                      ���������������``f� """""" ����f`������ ���������������                      ���������������ff``fj�� """ �����ff����� ���������������                      ���������������ffffff���� ������ff��������������������                      ��������������ff��`f���������  ��f`���������������������                      ��������������ff����hj�������n���ff���������������������                     ����� """"     fn�����`�������f����ff""   ����������������                     �����""""""""fn������`�����f�����f`"""""��������������                     ����"""""""""f�������f����fn�����f`""""" ���������������                     ����""""""""""f��������`���fn�����ff"""""����������������                    ���""""""""" ff���������`��f������ff"""""���������������                    ���"""""""""" ff���������fpfn������ff`"""""(���������������                    ��""""""""""" ff����������`�fn�����fff`""""""��������������                    �""""""""""" ff����������`�f������fff`""""""��������������                    �"""""""""""" ffn����������f������fff""""""(���������������                   """"""""""""*pffn����������f������fff"""""" ���������������                   """"""""""""�wff����������`f������ff`�"""""""��������������                   """""""""""�wwffn����������n�����fff`w�"""""""�������������                   """""""""(�www�fff���������������fff
ww"""""""(�������������                   """""""'�wwwwwpfffnn�������������ff`�ww�"""""""��������������                  """""""'wwwwwwwffff�������������ff`www�""""""" �������������                  """""""'zwwwwwwpffffn������������ff
www"""""""""�����������                  """""""'wwwwwwp�ffff������������ffwz""""""""""������������                  """"""""w�www�""��fffn�����������f`""""""""""""""(������������                 """"""""'wwz�""""w�fff����������ff`"""""""""""""""������������                 """""""""""""""""*��ffn����`f����ff"""""""""""""""(�����������                 """"""""""""""""""��ff����`fffffff""""""""""""""""����������                 """""""""""""""""""(�ffffff fffff`""""""""""""""""" ����������                 """"""""""""""""""""" fff`"""   """""""""""""""""""����������                """"""""""""""""""""""""""""""""""""""""""""""""""""" ����������                """"""""""""""""""""""""""""""""""""""""""""""""""""""���������                """""""""""""""""""""""""""""""""""""""""""""""""""""" ��������                                                                                                                                                                                                                ������������������������������������������                                     �������������������������������������������                                     ��������������������������������������������                                    ��������������������������������������������                                    �������������������� ���������������������                                    �����������������������������������������                                    ������������������������������������������                                    ���������������������������Ј����������������                                   ��������������������������������������������                                   ��������������������������������������������                                   ������������������ݍݍ������Ј���������������                                   ������������������ݍ������������������������                                  ������������������݌��ݍ���������������������                                  �����������������ݍ���ݍ���������������������                                  �����������������݈؍�ݍ�������������������                                  �����������������݆�`� ���݀����������������                                  �������������������f f�`���Ј����������������                                 ������������������� �������Ј����������������                                 ��������������������������������������� ������                                 �������������������������������������� ������                                 ������������������ؠn�f��f�������������������                                 �������������������n�Fn��f��������������������                                �������������������������f�����Ј��������������                                ���������������������N��f`������������������                                ������������������ݎ�L���f ���������������������                                �������������������������``������Ј��������������                               �������������������������`������Ј��������������                               ��������������������݀n`ff��������������������                               ����������������������ffnf������Ј������������                               ����������������������ff�f`������Ј�������������                               ����������������������nf���f2��������������������                              ������������������݈#&�����f#.���� ��������������                              ������������������n�rfn���n�#.��h��Ј�������������                              �������������������r�������'.������������������                              ��������������������r�������'r���Ј��������������                              ��������������������r�������'r���m����������������                             �������������������r�������'r���言      ��������                             �������������ݍ����2�������#r���h�����   �������                             �����������܌����3�������#r���`������  ��������                             ������������Ѐ����3.������#3.��`������  ���������                            �����������������3>������#3&�`������  ���������                            ����������������7r������7s n��������  ���������                            ������������������bww2&fn"7ww2n�������  ��������                            ������������������'wwwwwwwwwwrn�������� ���������                            ������������������'wwwwwwwwwww.�������� ����������                           ����������������n��7wwwwwwwwwww2�������� ����������                           ����������������n�#7wwwwwwwwwww2n�`������ ����������                           ������������������#7wwwwwwwwwww3.�`������ ���������                           ������������������37wwwwwwwwwwr3&�`�����������������                           ������������������33wwwww33www33 ������������������                          �����������������333ww33333w333&n������������������                          �����������������#3333333233332f` `����������������                          ���������������ffb333#7www2#3"
 n�������������������                          ���������������f�"33wwwww333 `��������������������                         ���������������fn�f337wwwwww33`��������������������                         ���������������fn��`337wwwwwws3`n��������������������                         ���������������fn��`""3wwwwwws3�������������������                         ���������������ff�f'ww"wwwws3"
�������������������                         ���������������ff`
���w�332'w� �`������������������                        ���������������n��������2z��p ���������������������                        ���������������n�`" ����*�p `���������������������                        ����������������n�f""  ���"""" n�����������������                        ����������������n��"""""
�""""" ��������������������                        ���������������n���""""""""""""" 0������� ��������������                       �������������������"""""""""""" 0������� ��������������                       ���������������n�f���""""""""" 3"������ �������������                       ����������������nn�  """""""" �f`������ �������������                       ������������������`""""""""" zfff������ ���������������                      ����������������f """"""""~��f`������ ���������������                      ���������������f f�� """""����f`������ ���������������                      ���������������ffffj��� ""�����ff��������������������                      ��������������ffffff���������ffff`���������������������                      ��������������fn����������n���f`����������������������                     �����   �����fn������������n���ff  �������������������                     �����"""""""" fn�����f������f�����f`"""""����������������                     �����"""""""""f�������`�����f�����f`"""""(��������������                     ����"""""""""f��������`����fn�����ff"""""���������������                     ����""""""""" ff�����������fn�����ff"""""���������������                    ���"""""""""" ff���������`wpff������ff"""""(���������������                    ��"""""""""" ff����������pfn������ff`""""" ��������������                    ��""""""""""" ff����������`�fn�����fff`""""""��������������                    �"""""""""""" ffn���������ff������fff`""""""��������������                    """"""""""""pffn����������f������fff"""""" ���������������                   """"""""""""'pffn����������`f������fff"""""""��������������                   """"""""""" �wff����������`n������ff`z""""""" �������������                   """"""""""(wwwffn���������������fff
wz"""""""�������������                   """""""*�wwwwwpfff�n�������������fffww�"""""" ��������������                  """""""'wwwwwwzffff�������������ff`�ww�"""""""(�������������                  """""""'zwwwwww�ffff�������������ff
www�""""""""������������                  """""""'zwwwwwwwfffn������������ff
wwz"""""""""(�����������                  """""""*w�wwwz""�fff������������f`" w�""""""""""������������                  """"""""�zwwx"""*zffn�����������f`"""""""""""""" ������������                 """"""""*w��"""""��ff������f����ff"""""""""""""""�����������                 """"""""""""""""""��fn����`fn��fff""""""""""""""" ����������                 """""""""""""""""" ��fffffffffff`"""""""""""""""""���������                 """""""""""""""""""" ffff`"" fff`""""""""""""""""" ����������                 """"""""""""""""""""""   """""""""""""""""""""""""""����������                """"""""""""""""""""""""""""""""""""""""""""""""""""" ����������                """"""""""""""""""""""""""""""""""""""""""""""""""""""��������                """""""""""""""""""""""""""""""""""""""""""""""""""""" ���������                                                                                                                                                                                                                